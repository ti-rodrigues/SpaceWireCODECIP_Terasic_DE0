// CPU.v

// Generated using ACDS version 13.1 162 at 2015.10.27.14:53:06

`timescale 1 ps / 1 ps
module CPU (
		input  wire        clk_clk,             //          clk.clk
		input  wire        reset_reset_n,       //        reset.reset_n
		output wire [11:0] sdram_addr,          //        sdram.addr
		output wire [1:0]  sdram_ba,            //             .ba
		output wire        sdram_cas_n,         //             .cas_n
		output wire        sdram_cke,           //             .cke
		output wire        sdram_cs_n,          //             .cs_n
		inout  wire [15:0] sdram_dq,            //             .dq
		output wire [1:0]  sdram_dqm,           //             .dqm
		output wire        sdram_ras_n,         //             .ras_n
		output wire        sdram_we_n,          //             .we_n
		output wire [6:0]  spw_tx_div_export,   //   spw_tx_div.export
		output wire [2:0]  spw_config_export,   //   spw_config.export
		output wire        spw_tick_in_export,  //  spw_tick_in.export
		output wire [7:0]  spw_time_in_export,  //  spw_time_in.export
		output wire        spw_reset_export,    //    spw_reset.export
		input  wire [2:0]  spw_state_export,    //    spw_state.export
		input  wire        spw_tick_o_export,   //   spw_tick_o.export
		input  wire [7:0]  spw_time_o_export,   //   spw_time_o.export
		input  wire [8:0]  spw_data_i_export,   //   spw_data_i.export
		input  wire        spw_tx_full_export,  //  spw_tx_full.export
		input  wire        spw_rx_empty_export, // spw_rx_empty.export
		output wire        spw_data_rd_export,  //  spw_data_rd.export
		output wire        spw_data_wr_export,  //  spw_data_wr.export
		output wire [8:0]  spw_data_o_export,   //   spw_data_o.export
		output wire [31:0] display7seg_export,  //  display7seg.export
		output wire [9:0]  led_export           //          led.export
	);

	wire   [1:0] mm_interconnect_0_spw_state_s1_address;                    // mm_interconnect_0:spw_state_s1_address -> spw_state:address
	wire  [31:0] mm_interconnect_0_spw_state_s1_readdata;                   // spw_state:readdata -> mm_interconnect_0:spw_state_s1_readdata
	wire   [1:0] mm_interconnect_0_spw_time_o_s1_address;                   // mm_interconnect_0:spw_time_o_s1_address -> spw_time_o:address
	wire  [31:0] mm_interconnect_0_spw_time_o_s1_readdata;                  // spw_time_o:readdata -> mm_interconnect_0:spw_time_o_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [24:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire   [1:0] mm_interconnect_0_spw_rx_empty_s1_address;                 // mm_interconnect_0:spw_rx_empty_s1_address -> spw_rx_empty:address
	wire  [31:0] mm_interconnect_0_spw_rx_empty_s1_readdata;                // spw_rx_empty:readdata -> mm_interconnect_0:spw_rx_empty_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_0_display7seg_s1_writedata;                // mm_interconnect_0:display7seg_s1_writedata -> display7seg:writedata
	wire   [1:0] mm_interconnect_0_display7seg_s1_address;                  // mm_interconnect_0:display7seg_s1_address -> display7seg:address
	wire         mm_interconnect_0_display7seg_s1_chipselect;               // mm_interconnect_0:display7seg_s1_chipselect -> display7seg:chipselect
	wire         mm_interconnect_0_display7seg_s1_write;                    // mm_interconnect_0:display7seg_s1_write -> display7seg:write_n
	wire  [31:0] mm_interconnect_0_display7seg_s1_readdata;                 // display7seg:readdata -> mm_interconnect_0:display7seg_s1_readdata
	wire  [31:0] mm_interconnect_0_spw_tx_div_s1_writedata;                 // mm_interconnect_0:spw_tx_div_s1_writedata -> spw_tx_div:writedata
	wire   [1:0] mm_interconnect_0_spw_tx_div_s1_address;                   // mm_interconnect_0:spw_tx_div_s1_address -> spw_tx_div:address
	wire         mm_interconnect_0_spw_tx_div_s1_chipselect;                // mm_interconnect_0:spw_tx_div_s1_chipselect -> spw_tx_div:chipselect
	wire         mm_interconnect_0_spw_tx_div_s1_write;                     // mm_interconnect_0:spw_tx_div_s1_write -> spw_tx_div:write_n
	wire  [31:0] mm_interconnect_0_spw_tx_div_s1_readdata;                  // spw_tx_div:readdata -> mm_interconnect_0:spw_tx_div_s1_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [24:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire  [31:0] mm_interconnect_0_spw_reset_s1_writedata;                  // mm_interconnect_0:spw_reset_s1_writedata -> spw_reset:writedata
	wire   [1:0] mm_interconnect_0_spw_reset_s1_address;                    // mm_interconnect_0:spw_reset_s1_address -> spw_reset:address
	wire         mm_interconnect_0_spw_reset_s1_chipselect;                 // mm_interconnect_0:spw_reset_s1_chipselect -> spw_reset:chipselect
	wire         mm_interconnect_0_spw_reset_s1_write;                      // mm_interconnect_0:spw_reset_s1_write -> spw_reset:write_n
	wire  [31:0] mm_interconnect_0_spw_reset_s1_readdata;                   // spw_reset:readdata -> mm_interconnect_0:spw_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_spw_data_i_s1_address;                   // mm_interconnect_0:spw_data_i_s1_address -> spw_data_i:address
	wire  [31:0] mm_interconnect_0_spw_data_i_s1_readdata;                  // spw_data_i:readdata -> mm_interconnect_0:spw_data_i_s1_readdata
	wire   [1:0] mm_interconnect_0_spw_tick_o_s1_address;                   // mm_interconnect_0:spw_tick_o_s1_address -> spw_tick_o:address
	wire  [31:0] mm_interconnect_0_spw_tick_o_s1_readdata;                  // spw_tick_o:readdata -> mm_interconnect_0:spw_tick_o_s1_readdata
	wire  [31:0] mm_interconnect_0_spw_tick_in_s1_writedata;                // mm_interconnect_0:spw_tick_in_s1_writedata -> spw_tick_in:writedata
	wire   [1:0] mm_interconnect_0_spw_tick_in_s1_address;                  // mm_interconnect_0:spw_tick_in_s1_address -> spw_tick_in:address
	wire         mm_interconnect_0_spw_tick_in_s1_chipselect;               // mm_interconnect_0:spw_tick_in_s1_chipselect -> spw_tick_in:chipselect
	wire         mm_interconnect_0_spw_tick_in_s1_write;                    // mm_interconnect_0:spw_tick_in_s1_write -> spw_tick_in:write_n
	wire  [31:0] mm_interconnect_0_spw_tick_in_s1_readdata;                 // spw_tick_in:readdata -> mm_interconnect_0:spw_tick_in_s1_readdata
	wire  [31:0] mm_interconnect_0_spw_data_rd_s1_writedata;                // mm_interconnect_0:spw_data_rd_s1_writedata -> spw_data_rd:writedata
	wire   [1:0] mm_interconnect_0_spw_data_rd_s1_address;                  // mm_interconnect_0:spw_data_rd_s1_address -> spw_data_rd:address
	wire         mm_interconnect_0_spw_data_rd_s1_chipselect;               // mm_interconnect_0:spw_data_rd_s1_chipselect -> spw_data_rd:chipselect
	wire         mm_interconnect_0_spw_data_rd_s1_write;                    // mm_interconnect_0:spw_data_rd_s1_write -> spw_data_rd:write_n
	wire  [31:0] mm_interconnect_0_spw_data_rd_s1_readdata;                 // spw_data_rd:readdata -> mm_interconnect_0:spw_data_rd_s1_readdata
	wire  [31:0] mm_interconnect_0_spw_time_in_s1_writedata;                // mm_interconnect_0:spw_time_in_s1_writedata -> spw_time_in:writedata
	wire   [1:0] mm_interconnect_0_spw_time_in_s1_address;                  // mm_interconnect_0:spw_time_in_s1_address -> spw_time_in:address
	wire         mm_interconnect_0_spw_time_in_s1_chipselect;               // mm_interconnect_0:spw_time_in_s1_chipselect -> spw_time_in:chipselect
	wire         mm_interconnect_0_spw_time_in_s1_write;                    // mm_interconnect_0:spw_time_in_s1_write -> spw_time_in:write_n
	wire  [31:0] mm_interconnect_0_spw_time_in_s1_readdata;                 // spw_time_in:readdata -> mm_interconnect_0:spw_time_in_s1_readdata
	wire  [31:0] mm_interconnect_0_spw_data_wr_s1_writedata;                // mm_interconnect_0:spw_data_wr_s1_writedata -> spw_data_wr:writedata
	wire   [1:0] mm_interconnect_0_spw_data_wr_s1_address;                  // mm_interconnect_0:spw_data_wr_s1_address -> spw_data_wr:address
	wire         mm_interconnect_0_spw_data_wr_s1_chipselect;               // mm_interconnect_0:spw_data_wr_s1_chipselect -> spw_data_wr:chipselect
	wire         mm_interconnect_0_spw_data_wr_s1_write;                    // mm_interconnect_0:spw_data_wr_s1_write -> spw_data_wr:write_n
	wire  [31:0] mm_interconnect_0_spw_data_wr_s1_readdata;                 // spw_data_wr:readdata -> mm_interconnect_0:spw_data_wr_s1_readdata
	wire  [31:0] mm_interconnect_0_spw_data_o_s1_writedata;                 // mm_interconnect_0:spw_data_o_s1_writedata -> spw_data_o:writedata
	wire   [1:0] mm_interconnect_0_spw_data_o_s1_address;                   // mm_interconnect_0:spw_data_o_s1_address -> spw_data_o:address
	wire         mm_interconnect_0_spw_data_o_s1_chipselect;                // mm_interconnect_0:spw_data_o_s1_chipselect -> spw_data_o:chipselect
	wire         mm_interconnect_0_spw_data_o_s1_write;                     // mm_interconnect_0:spw_data_o_s1_write -> spw_data_o:write_n
	wire  [31:0] mm_interconnect_0_spw_data_o_s1_readdata;                  // spw_data_o:readdata -> mm_interconnect_0:spw_data_o_s1_readdata
	wire   [1:0] mm_interconnect_0_spw_tx_full_s1_address;                  // mm_interconnect_0:spw_tx_full_s1_address -> spw_tx_full:address
	wire  [31:0] mm_interconnect_0_spw_tx_full_s1_readdata;                 // spw_tx_full:readdata -> mm_interconnect_0:spw_tx_full_s1_readdata
	wire  [31:0] mm_interconnect_0_spw_config_s1_writedata;                 // mm_interconnect_0:spw_config_s1_writedata -> spw_config:writedata
	wire   [1:0] mm_interconnect_0_spw_config_s1_address;                   // mm_interconnect_0:spw_config_s1_address -> spw_config:address
	wire         mm_interconnect_0_spw_config_s1_chipselect;                // mm_interconnect_0:spw_config_s1_chipselect -> spw_config:chipselect
	wire         mm_interconnect_0_spw_config_s1_write;                     // mm_interconnect_0:spw_config_s1_write -> spw_config:write_n
	wire  [31:0] mm_interconnect_0_spw_config_s1_readdata;                  // spw_config:readdata -> mm_interconnect_0:spw_config_s1_readdata
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire   [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu:reset_n, display7seg:reset_n, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset, sdram:reset_n, spw_config:reset_n, spw_data_i:reset_n, spw_data_o:reset_n, spw_data_rd:reset_n, spw_data_wr:reset_n, spw_reset:reset_n, spw_rx_empty:reset_n, spw_state:reset_n, spw_tick_in:reset_n, spw_tick_o:reset_n, spw_time_in:reset_n, spw_time_o:reset_n, spw_tx_div:reset_n, spw_tx_full:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]

	CPU_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                    //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	CPU_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	CPU_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)              //       .reset_req
	);

	CPU_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	CPU_spw_tx_div spw_tx_div (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_spw_tx_div_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_tx_div_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_tx_div_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_tx_div_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_tx_div_s1_readdata),   //                    .readdata
		.out_port   (spw_tx_div_export)                           // external_connection.export
	);

	CPU_spw_config spw_config (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_spw_config_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_config_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_config_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_config_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_config_s1_readdata),   //                    .readdata
		.out_port   (spw_config_export)                           // external_connection.export
	);

	CPU_spw_tick_in spw_tick_in (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_spw_tick_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_tick_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_tick_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_tick_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_tick_in_s1_readdata),   //                    .readdata
		.out_port   (spw_tick_in_export)                           // external_connection.export
	);

	CPU_spw_time_in spw_time_in (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_spw_time_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_time_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_time_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_time_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_time_in_s1_readdata),   //                    .readdata
		.out_port   (spw_time_in_export)                           // external_connection.export
	);

	CPU_spw_data_o spw_data_o (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_spw_data_o_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_data_o_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_data_o_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_data_o_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_data_o_s1_readdata),   //                    .readdata
		.out_port   (spw_data_o_export)                           // external_connection.export
	);

	CPU_spw_tick_in spw_data_wr (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_spw_data_wr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_data_wr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_data_wr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_data_wr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_data_wr_s1_readdata),   //                    .readdata
		.out_port   (spw_data_wr_export)                           // external_connection.export
	);

	CPU_spw_data_i spw_data_i (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_spw_data_i_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spw_data_i_s1_readdata), //                    .readdata
		.in_port  (spw_data_i_export)                         // external_connection.export
	);

	CPU_spw_tick_in spw_data_rd (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_spw_data_rd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_data_rd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_data_rd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_data_rd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_data_rd_s1_readdata),   //                    .readdata
		.out_port   (spw_data_rd_export)                           // external_connection.export
	);

	CPU_spw_rx_empty spw_rx_empty (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_spw_rx_empty_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spw_rx_empty_s1_readdata), //                    .readdata
		.in_port  (spw_rx_empty_export)                         // external_connection.export
	);

	CPU_spw_rx_empty spw_tx_full (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_spw_tx_full_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spw_tx_full_s1_readdata), //                    .readdata
		.in_port  (spw_tx_full_export)                         // external_connection.export
	);

	CPU_spw_time_o spw_time_o (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_spw_time_o_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spw_time_o_s1_readdata), //                    .readdata
		.in_port  (spw_time_o_export)                         // external_connection.export
	);

	CPU_spw_rx_empty spw_tick_o (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_spw_tick_o_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spw_tick_o_s1_readdata), //                    .readdata
		.in_port  (spw_tick_o_export)                         // external_connection.export
	);

	CPU_spw_state spw_state (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_spw_state_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spw_state_s1_readdata), //                    .readdata
		.in_port  (spw_state_export)                         // external_connection.export
	);

	CPU_spw_tick_in spw_reset (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_spw_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spw_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spw_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spw_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spw_reset_s1_readdata),   //                    .readdata
		.out_port   (spw_reset_export)                           // external_connection.export
	);

	CPU_display7seg display7seg (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_display7seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display7seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display7seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display7seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display7seg_s1_readdata),   //                    .readdata
		.out_port   (display7seg_export)                           // external_connection.export
	);

	CPU_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	CPU_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                                   //                         clk_0_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                   cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                  .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                  .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                  .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                  .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                  .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                  .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                  .readdata
		.cpu_jtag_debug_module_address           (mm_interconnect_0_cpu_jtag_debug_module_address),           //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write             (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                  .write
		.cpu_jtag_debug_module_read              (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                  .read
		.cpu_jtag_debug_module_readdata          (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                  .readdata
		.cpu_jtag_debug_module_writedata         (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                  .writedata
		.cpu_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                  .debugaccess
		.display7seg_s1_address                  (mm_interconnect_0_display7seg_s1_address),                  //                    display7seg_s1.address
		.display7seg_s1_write                    (mm_interconnect_0_display7seg_s1_write),                    //                                  .write
		.display7seg_s1_readdata                 (mm_interconnect_0_display7seg_s1_readdata),                 //                                  .readdata
		.display7seg_s1_writedata                (mm_interconnect_0_display7seg_s1_writedata),                //                                  .writedata
		.display7seg_s1_chipselect               (mm_interconnect_0_display7seg_s1_chipselect),               //                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.led_s1_address                          (mm_interconnect_0_led_s1_address),                          //                            led_s1.address
		.led_s1_write                            (mm_interconnect_0_led_s1_write),                            //                                  .write
		.led_s1_readdata                         (mm_interconnect_0_led_s1_readdata),                         //                                  .readdata
		.led_s1_writedata                        (mm_interconnect_0_led_s1_writedata),                        //                                  .writedata
		.led_s1_chipselect                       (mm_interconnect_0_led_s1_chipselect),                       //                                  .chipselect
		.onchip_memory2_s1_address               (mm_interconnect_0_onchip_memory2_s1_address),               //                 onchip_memory2_s1.address
		.onchip_memory2_s1_write                 (mm_interconnect_0_onchip_memory2_s1_write),                 //                                  .write
		.onchip_memory2_s1_readdata              (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                  .readdata
		.onchip_memory2_s1_writedata             (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                  .writedata
		.onchip_memory2_s1_byteenable            (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                  .byteenable
		.onchip_memory2_s1_chipselect            (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                  .chipselect
		.onchip_memory2_s1_clken                 (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                  .clken
		.sdram_s1_address                        (mm_interconnect_0_sdram_s1_address),                        //                          sdram_s1.address
		.sdram_s1_write                          (mm_interconnect_0_sdram_s1_write),                          //                                  .write
		.sdram_s1_read                           (mm_interconnect_0_sdram_s1_read),                           //                                  .read
		.sdram_s1_readdata                       (mm_interconnect_0_sdram_s1_readdata),                       //                                  .readdata
		.sdram_s1_writedata                      (mm_interconnect_0_sdram_s1_writedata),                      //                                  .writedata
		.sdram_s1_byteenable                     (mm_interconnect_0_sdram_s1_byteenable),                     //                                  .byteenable
		.sdram_s1_readdatavalid                  (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                  .readdatavalid
		.sdram_s1_waitrequest                    (mm_interconnect_0_sdram_s1_waitrequest),                    //                                  .waitrequest
		.sdram_s1_chipselect                     (mm_interconnect_0_sdram_s1_chipselect),                     //                                  .chipselect
		.spw_config_s1_address                   (mm_interconnect_0_spw_config_s1_address),                   //                     spw_config_s1.address
		.spw_config_s1_write                     (mm_interconnect_0_spw_config_s1_write),                     //                                  .write
		.spw_config_s1_readdata                  (mm_interconnect_0_spw_config_s1_readdata),                  //                                  .readdata
		.spw_config_s1_writedata                 (mm_interconnect_0_spw_config_s1_writedata),                 //                                  .writedata
		.spw_config_s1_chipselect                (mm_interconnect_0_spw_config_s1_chipselect),                //                                  .chipselect
		.spw_data_i_s1_address                   (mm_interconnect_0_spw_data_i_s1_address),                   //                     spw_data_i_s1.address
		.spw_data_i_s1_readdata                  (mm_interconnect_0_spw_data_i_s1_readdata),                  //                                  .readdata
		.spw_data_o_s1_address                   (mm_interconnect_0_spw_data_o_s1_address),                   //                     spw_data_o_s1.address
		.spw_data_o_s1_write                     (mm_interconnect_0_spw_data_o_s1_write),                     //                                  .write
		.spw_data_o_s1_readdata                  (mm_interconnect_0_spw_data_o_s1_readdata),                  //                                  .readdata
		.spw_data_o_s1_writedata                 (mm_interconnect_0_spw_data_o_s1_writedata),                 //                                  .writedata
		.spw_data_o_s1_chipselect                (mm_interconnect_0_spw_data_o_s1_chipselect),                //                                  .chipselect
		.spw_data_rd_s1_address                  (mm_interconnect_0_spw_data_rd_s1_address),                  //                    spw_data_rd_s1.address
		.spw_data_rd_s1_write                    (mm_interconnect_0_spw_data_rd_s1_write),                    //                                  .write
		.spw_data_rd_s1_readdata                 (mm_interconnect_0_spw_data_rd_s1_readdata),                 //                                  .readdata
		.spw_data_rd_s1_writedata                (mm_interconnect_0_spw_data_rd_s1_writedata),                //                                  .writedata
		.spw_data_rd_s1_chipselect               (mm_interconnect_0_spw_data_rd_s1_chipselect),               //                                  .chipselect
		.spw_data_wr_s1_address                  (mm_interconnect_0_spw_data_wr_s1_address),                  //                    spw_data_wr_s1.address
		.spw_data_wr_s1_write                    (mm_interconnect_0_spw_data_wr_s1_write),                    //                                  .write
		.spw_data_wr_s1_readdata                 (mm_interconnect_0_spw_data_wr_s1_readdata),                 //                                  .readdata
		.spw_data_wr_s1_writedata                (mm_interconnect_0_spw_data_wr_s1_writedata),                //                                  .writedata
		.spw_data_wr_s1_chipselect               (mm_interconnect_0_spw_data_wr_s1_chipselect),               //                                  .chipselect
		.spw_reset_s1_address                    (mm_interconnect_0_spw_reset_s1_address),                    //                      spw_reset_s1.address
		.spw_reset_s1_write                      (mm_interconnect_0_spw_reset_s1_write),                      //                                  .write
		.spw_reset_s1_readdata                   (mm_interconnect_0_spw_reset_s1_readdata),                   //                                  .readdata
		.spw_reset_s1_writedata                  (mm_interconnect_0_spw_reset_s1_writedata),                  //                                  .writedata
		.spw_reset_s1_chipselect                 (mm_interconnect_0_spw_reset_s1_chipselect),                 //                                  .chipselect
		.spw_rx_empty_s1_address                 (mm_interconnect_0_spw_rx_empty_s1_address),                 //                   spw_rx_empty_s1.address
		.spw_rx_empty_s1_readdata                (mm_interconnect_0_spw_rx_empty_s1_readdata),                //                                  .readdata
		.spw_state_s1_address                    (mm_interconnect_0_spw_state_s1_address),                    //                      spw_state_s1.address
		.spw_state_s1_readdata                   (mm_interconnect_0_spw_state_s1_readdata),                   //                                  .readdata
		.spw_tick_in_s1_address                  (mm_interconnect_0_spw_tick_in_s1_address),                  //                    spw_tick_in_s1.address
		.spw_tick_in_s1_write                    (mm_interconnect_0_spw_tick_in_s1_write),                    //                                  .write
		.spw_tick_in_s1_readdata                 (mm_interconnect_0_spw_tick_in_s1_readdata),                 //                                  .readdata
		.spw_tick_in_s1_writedata                (mm_interconnect_0_spw_tick_in_s1_writedata),                //                                  .writedata
		.spw_tick_in_s1_chipselect               (mm_interconnect_0_spw_tick_in_s1_chipselect),               //                                  .chipselect
		.spw_tick_o_s1_address                   (mm_interconnect_0_spw_tick_o_s1_address),                   //                     spw_tick_o_s1.address
		.spw_tick_o_s1_readdata                  (mm_interconnect_0_spw_tick_o_s1_readdata),                  //                                  .readdata
		.spw_time_in_s1_address                  (mm_interconnect_0_spw_time_in_s1_address),                  //                    spw_time_in_s1.address
		.spw_time_in_s1_write                    (mm_interconnect_0_spw_time_in_s1_write),                    //                                  .write
		.spw_time_in_s1_readdata                 (mm_interconnect_0_spw_time_in_s1_readdata),                 //                                  .readdata
		.spw_time_in_s1_writedata                (mm_interconnect_0_spw_time_in_s1_writedata),                //                                  .writedata
		.spw_time_in_s1_chipselect               (mm_interconnect_0_spw_time_in_s1_chipselect),               //                                  .chipselect
		.spw_time_o_s1_address                   (mm_interconnect_0_spw_time_o_s1_address),                   //                     spw_time_o_s1.address
		.spw_time_o_s1_readdata                  (mm_interconnect_0_spw_time_o_s1_readdata),                  //                                  .readdata
		.spw_tx_div_s1_address                   (mm_interconnect_0_spw_tx_div_s1_address),                   //                     spw_tx_div_s1.address
		.spw_tx_div_s1_write                     (mm_interconnect_0_spw_tx_div_s1_write),                     //                                  .write
		.spw_tx_div_s1_readdata                  (mm_interconnect_0_spw_tx_div_s1_readdata),                  //                                  .readdata
		.spw_tx_div_s1_writedata                 (mm_interconnect_0_spw_tx_div_s1_writedata),                 //                                  .writedata
		.spw_tx_div_s1_chipselect                (mm_interconnect_0_spw_tx_div_s1_chipselect),                //                                  .chipselect
		.spw_tx_full_s1_address                  (mm_interconnect_0_spw_tx_full_s1_address),                  //                    spw_tx_full_s1.address
		.spw_tx_full_s1_readdata                 (mm_interconnect_0_spw_tx_full_s1_readdata)                  //                                  .readdata
	);

	CPU_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
